module inst_mem #(
    parameter inst_SIZE =   16,
    parameter PC_SIZE   =   13
) (
    input   wire    [PC_SIZE-1:0]       PC,

    output  wire    [inst_SIZE-1:0]     instruction
);
    


endmodule