module MUX_2_to_1 (
    ports
);
    
endmodule