module ALU #(
    parameter inst_SIZE = 16
) (
    input   wire    [2:0]               alu_ctrl,
    input   wire    [inst_SIZE-1:0]     read_data_1,
    input   wire    [inst_SIZE-1:0]     read_data_2,

    output  wire                        zero,
    output          
);
    
endmodule