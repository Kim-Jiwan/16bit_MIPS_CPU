module moduleName #(
    parameter inst_SIZE = 16
) (
    input   wire                        PC,

    output  wire    [inst_SIZE-1:0]     instruction
);
    


endmodule