module ALU (
    input   wire    [2:0]   alu_ctrl,
    input   wire    [15:0]  read_data_1,
    input   wire    [15:0]  read_data_2,

    output  wire            zero,
    output          
);
    
endmodule