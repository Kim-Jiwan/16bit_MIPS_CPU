module cpu (
    input   wire    clk,
    input   wire    rst
);
    
endmodule